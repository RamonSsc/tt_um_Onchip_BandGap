VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Onchip_BandGap
  CLASS BLOCK ;
  FOREIGN tt_um_Onchip_BandGap ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.422000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 50.000000 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 6.750000 ;
    ANTENNADIFFAREA 0.148500 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VSS
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 457.036774 ;
    PORT
      LAYER met4 ;
        RECT 30.000 5.000 35.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.000 5.000 55.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.000 5.000 115.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.000 5.000 75.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.000 5.000 95.000 220.760 ;
    END
  END VSS
  PIN VDPWR
    PORT
      LAYER met4 ;
        RECT 20.000 5.000 25.000 220.760 ;
    END
  END VDPWR
  PIN VDD
    ANTENNAGATEAREA 514.519958 ;
    ANTENNADIFFAREA 510.403992 ;
    PORT
      LAYER met4 ;
        RECT 80.000 5.000 85.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.000 5.000 45.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.000 5.000 65.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.000 5.000 105.000 220.760 ;
    END
  END VDD
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 10.000 5.000 15.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 36.540 34.560 111.520 202.935 ;
      LAYER li1 ;
        RECT 36.850 34.690 111.210 202.805 ;
      LAYER met1 ;
        RECT 30.000 32.665 124.815 206.415 ;
      LAYER met2 ;
        RECT 30.000 32.665 124.815 206.415 ;
      LAYER met3 ;
        RECT 30.000 34.690 154.260 206.415 ;
      LAYER met4 ;
        RECT 10.000 224.360 30.270 224.760 ;
        RECT 31.370 224.360 33.030 224.760 ;
        RECT 34.130 224.360 35.790 224.760 ;
        RECT 36.890 224.360 38.550 224.760 ;
        RECT 39.650 224.360 41.310 224.760 ;
        RECT 42.410 224.360 44.070 224.760 ;
        RECT 45.170 224.360 46.830 224.760 ;
        RECT 47.930 224.360 49.590 224.760 ;
        RECT 50.690 224.360 52.350 224.760 ;
        RECT 53.450 224.360 55.110 224.760 ;
        RECT 56.210 224.360 57.870 224.760 ;
        RECT 58.970 224.360 60.630 224.760 ;
        RECT 61.730 224.360 63.390 224.760 ;
        RECT 64.490 224.360 66.150 224.760 ;
        RECT 67.250 224.360 68.910 224.760 ;
        RECT 70.010 224.360 71.670 224.760 ;
        RECT 72.770 224.360 74.430 224.760 ;
        RECT 75.530 224.360 77.190 224.760 ;
        RECT 78.290 224.360 79.950 224.760 ;
        RECT 81.050 224.360 82.710 224.760 ;
        RECT 83.810 224.360 85.470 224.760 ;
        RECT 86.570 224.360 88.230 224.760 ;
        RECT 89.330 224.360 90.990 224.760 ;
        RECT 92.090 224.360 93.750 224.760 ;
        RECT 94.850 224.360 96.510 224.760 ;
        RECT 97.610 224.360 99.270 224.760 ;
        RECT 100.370 224.360 102.030 224.760 ;
        RECT 103.130 224.360 104.790 224.760 ;
        RECT 105.890 224.360 107.550 224.760 ;
        RECT 108.650 224.360 110.310 224.760 ;
        RECT 111.410 224.360 113.070 224.760 ;
        RECT 114.170 224.360 115.830 224.760 ;
        RECT 116.930 224.360 118.590 224.760 ;
        RECT 119.690 224.360 121.350 224.760 ;
        RECT 122.450 224.360 124.110 224.760 ;
        RECT 125.210 224.360 126.870 224.760 ;
        RECT 127.970 224.360 129.630 224.760 ;
        RECT 130.730 224.360 132.390 224.760 ;
        RECT 133.490 224.360 135.150 224.760 ;
        RECT 136.250 224.360 137.910 224.760 ;
        RECT 139.010 224.360 140.670 224.760 ;
        RECT 141.770 224.360 143.430 224.760 ;
        RECT 144.530 224.360 146.190 224.760 ;
        RECT 147.290 224.360 154.260 224.760 ;
        RECT 10.000 221.160 154.260 224.360 ;
        RECT 10.000 220.760 15.000 221.160 ;
        RECT 15.400 4.600 19.600 221.160 ;
        RECT 25.400 4.600 29.600 221.160 ;
        RECT 35.400 4.600 39.600 221.160 ;
        RECT 45.400 4.600 49.600 221.160 ;
        RECT 55.400 4.600 59.600 221.160 ;
        RECT 65.400 4.600 69.600 221.160 ;
        RECT 75.400 4.600 79.600 221.160 ;
        RECT 85.400 4.600 89.600 221.160 ;
        RECT 95.400 4.600 99.600 221.160 ;
        RECT 105.400 4.600 109.600 221.160 ;
        RECT 115.400 4.600 154.260 221.160 ;
        RECT 10.000 1.400 154.260 4.600 ;
        RECT 10.000 1.000 16.170 1.400 ;
        RECT 17.870 1.000 35.490 1.400 ;
        RECT 37.190 1.000 54.810 1.400 ;
        RECT 56.510 1.000 74.130 1.400 ;
        RECT 75.830 1.000 93.450 1.400 ;
        RECT 95.150 1.000 112.770 1.400 ;
        RECT 114.470 1.000 132.090 1.400 ;
        RECT 133.790 1.000 151.410 1.400 ;
        RECT 153.110 1.000 154.260 1.400 ;
  END
END tt_um_Onchip_BandGap
END LIBRARY

